module ram();

parameter size = 256; //256 line * 4 bytes/line

reg [31:0] ram [size-1:0] // memory matrix, unit in words 

endmodule


