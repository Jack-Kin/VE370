module 2way_wb();



endmodule
