module 2way_wt();


endmodule
